/**************************
          control
***************************/

`define USE_SWITCH
//`define COMPILE_FRAME
`define COMPILE_SMALL

/**************************
          color
***************************/

//background
`define STATUS_BAR_COLOR  24'h7f7f7f
`define GROUND_COLOR  24'hffffff

//shell
`define SHELL_0 24'hff0000
`define SHELL_1 24'h0000ff

//wall
`define WALL_0 24'hffff00
`define WALL_1 24'h00ffff