/**************************
          control
***************************/

`define USE_SWITCH
//`define COMPILE_FRAME
`define COMPILE_SMALL
`define COMPILE_MULTIPLE_MAPS

/**************************
          color
***************************/

//background
`define STATUS_BAR_COLOR  24'hadadad
`define GROUND_COLOR  24'hffffff

//shell
`define SHELL_0 24'hff0000
`define SHELL_1 24'h0000ff

//wall
`define WALL_0 24'h548c00
`define WALL_1 24'h00ec00
`define WALL_2 24'h02df82
`define WALL_3 24'h8cea00

//life
`define TANK_LIFE 5
`define WALL_LIFE 3