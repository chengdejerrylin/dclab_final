//control
//`define COMPILE_FRAME

//color
`define STATUS_BAR_COLOR  24'h7f7f7f
`define GROUND_COLOR  24'h00ff00