`define COMPILE_FRAME